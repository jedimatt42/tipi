`ifndef _shift_pload_sout_vh_
`define _shift_pload_sout_vh_

module shift_pload_sout (
    // Clock for shifting
    input clk,
	 // Select
	 input select,
	 // load tmp with data to shift out.
    input aload,
	 // Data to load from
    input [7:0]data,
	 // output bit from the left.
    output sout
);

reg [7:0]tmp;

always @(posedge clk) begin
  if (aload && select) tmp = data;
  else if (select) tmp = { tmp[6:0], 1'b0 };
end

assign sout = tmp[7];

endmodule

`endif
